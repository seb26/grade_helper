<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>seb_bimok_apple_bnw_tinted</Description>
				<Slope>1.00000 1.00000 1.00000</Slope>
				<Offset>0.00000 0.00000 0.00000</Offset>
				<Power>1.00000 1.00000 1.00000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
