<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A014C004_220609_R111">
			<SOPNode>
				<Slope>0.700893 0.673690 0.649528</Slope>
				<Offset>0.002119 -0.006529 -0.027731</Offset>
				<Power>0.963005 0.952813 1.002028</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
