<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rr (modified)</Description>
				<Slope>0.74598 0.71701 0.69204</Slope>
				<Offset>0.00906 -0.00033 -0.02341</Offset>
				<Power>1.00509 0.99350 1.04940</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
