<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rrr (modified)</Description>
				<Slope>0.75131 0.72234 0.69737</Slope>
				<Offset>0.01275 0.00336 -0.01972</Offset>
				<Power>1.02724 1.01564 1.07154</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
