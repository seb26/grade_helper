<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description></Description>
				<Slope>1.22191 1.11508 1.08196</Slope>
				<Offset>-0.04047 0.00953 0.02475</Offset>
				<Power>1.00000 1.00000 1.00000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
