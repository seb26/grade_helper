<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description></Description>
				<Slope>0.96100 1.00439 1.07132</Slope>
				<Offset>-0.01588 0.00770 -0.02954</Offset>
				<Power>0.96739 1.01553 0.94217</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
