<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rrr (modified)</Description>
				<Slope>0.70745 0.67847 0.65351</Slope>
				<Offset>0.01275 0.00336 -0.01972</Offset>
				<Power>1.11713 1.10553 1.16143</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
