<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>New Look 1 (modified)</Description>
				<Slope>1.04785 0.98530 0.98793</Slope>
				<Offset>0.05747 0.00770 -0.08532</Offset>
				<Power>0.88370 1.03276 1.02384</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
