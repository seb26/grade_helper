<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rr (modified)</Description>
				<Slope>0.80167 0.77270 0.74773</Slope>
				<Offset>-0.01879 -0.02818 -0.05126</Offset>
				<Power>1.00509 0.99350 1.04940</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
