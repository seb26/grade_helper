<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description></Description>
				<Slope>1.08651 0.97968 0.94656</Slope>
				<Offset>-0.04047 0.00953 0.02475</Offset>
				<Power>1.00000 1.00000 1.00000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
