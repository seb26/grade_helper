<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description></Description>
				<Slope>1.0904 0.9810 0.9222</Slope>
				<Offset>0.0734 0.0000 -0.0558</Offset>
				<Power>0.9135 1.0170 1.0867</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
