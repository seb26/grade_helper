<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>emb_seb_v1_xx (modified) 4 (modified)</Description>
				<Slope>0.78851 0.78851 0.78851</Slope>
				<Offset>0.01123 -0.00234 -0.01720</Offset>
				<Power>1.00000 1.00000 1.00000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
