<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rrr</Description>
				<Slope>0.77856 0.74959 0.72462</Slope>
				<Offset>0.00160 -0.01370 -0.02560</Offset>
				<Power>0.95037 0.93877 0.99467</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
