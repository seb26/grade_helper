<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="cdl 3+4 lattice">
			<SOPNode>
				<Slope>0.853270 0.785874 0.772013</Slope>
				<Offset>0.056846 0.004464 -0.085888</Offset>
				<Power>0.791110 0.943110 0.958890</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
