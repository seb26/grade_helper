<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>rr</Description>
				<Slope>0.75889 0.72992 0.70496</Slope>
				<Offset>0.00906 -0.00033 -0.02341</Offset>
				<Power>1.00509 0.99350 1.04940</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
