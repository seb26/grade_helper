<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A009C008_220320_R4DG">
			<SOPNode>
				<Slope>0.928000 0.939958 0.951445</Slope>
				<Offset>-0.004923 -0.004987 -0.005047</Offset>
				<Power>1.000000 1.000000 1.000000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
