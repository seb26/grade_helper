<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A013C001_220609_R111">
			<SOPNode>
				<Slope>0.851631 0.851406 0.851159</Slope>
				<Offset>0.013529 0.000004 -0.014798</Offset>
				<Power>0.914900 0.914130 0.907720</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
