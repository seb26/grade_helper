<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A012C002_220609_R111">
			<SOPNode>
				<Slope>0.797080 0.797080 0.797080</Slope>
				<Offset>0.011760 -0.001810 -0.016670</Offset>
				<Power>0.915100 0.915100 0.915100</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
