<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A012C004_220609_R111">
			<SOPNode>
				<Slope>0.755136 0.753406 0.751522</Slope>
				<Offset>-0.038319 -0.049908 -0.062537</Offset>
				<Power>0.717036 0.716433 0.711409</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
