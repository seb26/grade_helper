<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>New Look 1 (modified)</Description>
				<Slope>0.83524 0.78538 0.78748</Slope>
				<Offset>0.06927 0.00590 -0.10202</Offset>
				<Power>0.80867 0.94508 0.93692</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
