<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A016C003_220609_R111">
			<SOPNode>
				<Slope>1.000000 1.000000 1.000000</Slope>
				<Offset>0.000000 0.000000 0.000000</Offset>
				<Power>1.000000 1.000000 1.000000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
