<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A006C005_220319_R4DG">
			<SOPNode>
				<Slope>1.230066 1.230066 1.230066</Slope>
				<Offset>-0.072518 -0.072518 -0.072518</Offset>
				<Power>0.834144 0.834144 0.834144</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
