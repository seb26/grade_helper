<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection>
			<SOPNode>
				<Description>emb_seb_v1_xx (modified) 4 (modified)</Description>
				<Slope>0.92019 0.92019 0.92019</Slope>
				<Offset>0.01176 -0.00181 -0.01667</Offset>
				<Power>0.91510 0.91510 0.91510</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.00000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
