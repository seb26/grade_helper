<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="A001C001_220319_R4DG">
			<SOPNode>
				<Slope>1.039667 1.039667 1.039667</Slope>
				<Offset>-0.060561 -0.060561 -0.060561</Offset>
				<Power>1.000000 1.000000 1.000000</Power>
			</SOPNode>
			<SATNode>
				<Saturation>1.000000</Saturation>
			</SATNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
